module round (
	input [31:0] first_32_bit,
	input [31:0] second_32_bit,
	input [127:0] sum,
	output [31:0] first_32_bit,
	output [31:0] second_32_bit
);

	


endmodule
