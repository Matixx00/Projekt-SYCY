/*
 * by SYCY_Proj_3
 *
 * Scheduler for several parallel synchronized TEA decryptors
 *
 *
 */
 
module input_scheduler (
	input			clk, rst,
			[63:0] 	in_word64,
			
	output	[63:0]	out_word64
	
);

endmodule
