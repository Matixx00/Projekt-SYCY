module miktea ();
endmodule
